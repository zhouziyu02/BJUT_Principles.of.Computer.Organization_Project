library verilog;
use verilog.vl_types.all;
entity ALU is
    port(
        A               : in     vl_logic_vector(31 downto 0);
        B               : in     vl_logic_vector(31 downto 0);
        ALU_op          : in     vl_logic_vector(2 downto 0);
        zero            : out    vl_logic;
        alu_out         : out    vl_logic_vector(31 downto 0);
        overflow        : out    vl_logic;
        slt             : in     vl_logic;
        addi            : in     vl_logic
    );
end ALU;
